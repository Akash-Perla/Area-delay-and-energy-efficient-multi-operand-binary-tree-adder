module BTA_CLA_tb#(parameter N=8,m=16);
reg clk;
reg [m-1:0]A,B,C,D,E,F,G,H;
reg C0;
wire [m+2:0]sum;
wire carry;

BTA_CLA_8 a1(clk,A,B,C,D,E,F,G,H,C0,sum,carry);

//initial repeat(255) #10 {A,B} = {A,B} + 8'b1;


initial begin

$dumpfile("BTA_CLA.vcd");
$dumpvars(0,BTA_CLA_tb);
end

initial begin
clk=0;
A=16'b0; B=16'b0; C=16'b0;D=16'b0;E=16'b0;F=16'b0;G=16'B0;H=16'b0; C0=0;
#20 A=16'b0101111000111010; B=16'b1111000010101110;C=16'b0101101011001010; D=16'b0110101100111110;E=16'b0101100100111010; F=16'b0100100000001110;G=16'b0011100111011010; H=16'b0101110010111110;
#20 A=16'b111001100001111; B=16'b0000010010111111;C=16'b0110100101111011; D=16'b0000100000011000;E=16'b1111010111000111; F=16'b0101100001000110;G=16'b0001001000111001; H=16'b0101001110101111;
//#20 A=16'b1110111010101101; B=16'b0010101001101110;
//#20 A=16'b1101010111011011; B=16'b1111111111111111;
#100 $finish;

end
always begin
#1 clk=~clk;
end

endmodule
